library verilog;
use verilog.vl_types.all;
entity tb_ifc_sv_unit is
end tb_ifc_sv_unit;
