/***********************************************************************
 * A SystemVerilog testbench for an instruction register; This file
 * contains the interface to connect the testbench to the design
 **********************************************************************/
 import instr_register_pkg::*;
interface tb_ifc (input logic clk);
 // timeunit 1ns/1ns;
 logic          load_en;
 logic          reset_n;
 opcode_t       opcode;
 operand_t      operand_a, operand_b;
 operand_t      result;
 address_t      write_pointer, read_pointer;
 instruction_t  instruction_word;


 clocking cb @(clk);
    output load_en;
    output reset_n;
    output opcode;
    output operand_a;
    output operand_b;
    output write_pointer;
    output read_pointer;
	  input result;
    input instruction_word;
 endclocking
 modport  TEST (clocking cb
 ); 
 

  // user-defined types are defined in instr_register_pkg.sv
  


  // ADD CODE TO DECLARE THE INTERFACE SIGNALS


endinterface: tb_ifc

